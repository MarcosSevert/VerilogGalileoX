`timescale 1ns/10ps

module demux_TB();
  reg in;
  reg [1:0] select;
  wire out3, out2, out1, out0;

  Demux_1_4 my_demux(in,select,{out3,out2,out1,out0});
  always #3 in=~in;

  initial begin
    $dumpfile("out.vcd");
    $dumpvars(1,demux_TB);
    in=0;

    select=2'b00;
    #20
    select=2'b01;
    #20
    select=2'b10;
    #20
    select=2'b11;
    #20
    $finish;
  end
  endmodule
